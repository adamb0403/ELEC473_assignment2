library verilog;
use verilog.vl_types.all;
entity tx_single_pulser_vlg_vec_tst is
end tx_single_pulser_vlg_vec_tst;
