library verilog;
use verilog.vl_types.all;
entity rx_shift_register_vlg_vec_tst is
end rx_shift_register_vlg_vec_tst;
