library verilog;
use verilog.vl_types.all;
entity irda_encoder_vlg_vec_tst is
end irda_encoder_vlg_vec_tst;
