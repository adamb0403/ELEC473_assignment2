library verilog;
use verilog.vl_types.all;
entity tx_shift_register_vlg_vec_tst is
end tx_shift_register_vlg_vec_tst;
