library verilog;
use verilog.vl_types.all;
entity tx_uart_vlg_vec_tst is
end tx_uart_vlg_vec_tst;
