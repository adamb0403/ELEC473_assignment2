library verilog;
use verilog.vl_types.all;
entity full_uart_vlg_vec_tst is
end full_uart_vlg_vec_tst;
