library verilog;
use verilog.vl_types.all;
entity irda_inverter_vlg_vec_tst is
end irda_inverter_vlg_vec_tst;
