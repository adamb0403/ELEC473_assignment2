library verilog;
use verilog.vl_types.all;
entity tx_baud_counter_vlg_vec_tst is
end tx_baud_counter_vlg_vec_tst;
