library verilog;
use verilog.vl_types.all;
entity tx_7segdecoder_vlg_vec_tst is
end tx_7segdecoder_vlg_vec_tst;
