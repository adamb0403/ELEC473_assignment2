library verilog;
use verilog.vl_types.all;
entity tx_controller_vlg_vec_tst is
end tx_controller_vlg_vec_tst;
