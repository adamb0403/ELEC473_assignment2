library verilog;
use verilog.vl_types.all;
entity rx_controller_vlg_vec_tst is
end rx_controller_vlg_vec_tst;
