library verilog;
use verilog.vl_types.all;
entity tx_parity_vlg_vec_tst is
end tx_parity_vlg_vec_tst;
