library verilog;
use verilog.vl_types.all;
entity tx_synchroniser_vlg_vec_tst is
end tx_synchroniser_vlg_vec_tst;
