library verilog;
use verilog.vl_types.all;
entity rx_parity_check_vlg_vec_tst is
end rx_parity_check_vlg_vec_tst;
